module top(...);
    input clk;
    output [3:0] led;

endmodule
